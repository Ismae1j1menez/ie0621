

`include "scoreboard.sv"
`include "stimulus.sv"
`include "monitor.sv"

`include "driver_bus_master.sv"
`include "interface_bus_master.sv"
`include "env.sv"
`include "tb_top.sv"
`include "test1.sv"
//`include "test2.sv"
//`include "test3.sv"
`include "mt48lc8m8a2.v"


