`include "top_hvl.sv"
`include "interface_bus_master.sv"
`include "driver.sv"
`include "scoreboard.sv"
`include "monitor.sv"
`include "agent.sv"
`include "env.sv"
`include "test_1.sv"
//`include "IS42VM16400K.V"
`include "mt48lc8m8a2.v"
`include "mt48lc2m32b2.v"