`include "IS42VM16400K.V"
`include "mt48lc8m8a2.v"
`include "mt48lc2m32b2.v"
