/********************************************************************
*  General Code Description
*  This code implements three important elements in a UVM verification 
*  environment: the `item`, the `sequences`, and the `driver`.
*  - `sdram_item`: Represents a transactional element with several 
*    properties that can be randomized.
*  - `gen_item_seq`: Generates a sequence of `sdram_item` elements to be 
*    processed.
*  - `sdram_driver`: Controls the bus and SDRAM interface, executing 
*    read and write operations based on the items generated by the sequence.
********************************************************************/

//------------------------------------------------------------------
// `sdram_item` Class
// Represents a transactional element in a UVM sequence, with 
// several fields that can be randomized and used in bus operations 
// (read/write).
//------------------------------------------------------------------
class sdram_item extends uvm_sequence_item;

  // UVM macros for automating the creation of methods and registering fields.
  `uvm_object_utils_begin(sdram_item)
  `uvm_field_int(writte, UVM_ALL_ON)     
  `uvm_field_int(bl, UVM_ALL_ON)         
  `uvm_field_int(amount_times, UVM_ALL_ON)
  `uvm_field_int(Address, UVM_ALL_ON)    
  `uvm_field_int(command, UVM_ALL_ON)    
  `uvm_field_int(delay, UVM_ALL_ON)      
  `uvm_field_int(iterations, UVM_ALL_ON) 
  `uvm_field_int(iteration_write, UVM_ALL_ON)
  `uvm_field_int(iteration_read, UVM_ALL_ON)
  `uvm_object_utils_end

  // Constructor to initialize the name of the sequence item.
  function new(string name = "sdram_item");
    super.new(name);
  endfunction

  // Declaration of random variables for the transaction.
  randc bit [31:0] writte;
  rand bit [7:0] bl;
  randc bit [7:0] amount_times;
  rand bit [31:0] Address;
  rand bit [1:0] command;
  rand bit [7:0] delay;
  rand bit [3:0] iterations;
  rand bit [2:0] iteration_write;
  rand bit [2:0] iteration_read;

  // Constraints to ensure valid values during simulation.
  constraint bl_c { bl >= 8 && bl <= 15; } 
  constraint amount_times_c { amount_times inside {[1:255]}; } 
  constraint command_c { command inside {0, 1}; } 
  constraint delay_c { delay inside {[1:255]}; } 
  constraint iterations_c { iterations inside {1, 2, 3, 4}; } 
  constraint address_c { Address inside {[32'h00000000 : 32'h00000FFC]}; } 
  
endclass


//------------------------------------------------------------------
// `gen_item_seq` Class
// Generates a sequence of `sdram_item` elements to be processed 
// in the UVM simulation.
//------------------------------------------------------------------
class gen_item_seq extends uvm_sequence #(sdram_item);

  // UVM macro to facilitate the creation and registration of the sequence.
  `uvm_object_utils(gen_item_seq)

  // Constructor to initialize an instance of the sequence.
  function new(string name="gen_item_seq");
    super.new(name);
  endfunction

  // Random variable that determines the number of items to generate.
  rand int num;
  
  // Constraint to ensure that the number of items is between 2 and 5.
  constraint c1 { num inside {[2:5]}; }

  // The body of the sequence that generates the `sdram_item` elements.
  virtual task body();
    for (int i = 0; i < num; i++) begin
      sdram_item f_item = sdram_item::type_id::create("f_item"); // Create a new item.

      start_item(f_item);          // Start the transaction.
      f_item.randomize();          // Randomize the fields of the item.
      `uvm_info("SEQ", $sformatf("Generate new item: command = %0d, address = %h", f_item.command, f_item.Address), UVM_LOW)
      f_item.print();              // Print the details of the generated item.
      finish_item(f_item);         // Finish the transaction.
    end
    `uvm_info("SEQ", $sformatf("Done generation of %0d items", num), UVM_LOW)
  endtask
endclass


//------------------------------------------------------------------
// `sdram_driver` Class
// Controls the bus and SDRAM interface, executing read and write 
// operations based on the items generated by the `gen_item_seq` sequence.
//------------------------------------------------------------------
class sdram_driver extends uvm_driver #(sdram_item);
  
  `uvm_component_utils(sdram_driver) // Macro to register the component in UVM.

  uvm_analysis_port #(sdram_item) analysis_port; // Analysis port to transmit transactions.

  // Constructor to initialize the driver.
  function new (string name = "sdram_driver", uvm_component parent = null);
    super.new(name, parent);
    analysis_port = new("analysis_port", this); // Initialize the analysis port.
  endfunction

  virtual interface_bus_master vif; // Virtual interface 

  // Build phase method to retrieve the virtual interface.
  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    if (!uvm_config_db #(virtual interface_bus_master)::get(this, "", "VIRTUAL_INTERFACE", vif)) begin
      `uvm_fatal("INTERFACE_CONNECT", "Failed to obtain virtual interface for the testbench")
    end
  endfunction

  // Connect phase method.
  virtual function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
  endfunction

  // Main run phase method for the driver, which handles the transactions.
  virtual task run_phase(uvm_phase phase);
    super.run_phase(phase);
    forever begin
      sdram_item f_item; 
      `uvm_info("DRV", $sformatf("Waiting for item from sequencer"), UVM_LOW)
      seq_item_port.get_next_item(f_item);

      if (f_item.command == 0) begin
        burst_write(f_item);
      end else if (f_item.command == 1) begin
        burst_read(f_item.Address);
      end

      analysis_port.write(f_item); 
      seq_item_port.item_done(); 
    end
  endtask

  // Reset task to initialize and reset signals.
  virtual task reset();
    vif.wb_addr_i      = 0;
    vif.wb_dat_i       = 0;
    vif.wb_sel_i       = 4'h0;
    vif.wb_we_i        = 1;
    vif.wb_stb_i       = 0;
    vif.wb_cyc_i       = 0;
    vif.RESETN         = 1'h1;
    #100

    vif.RESETN         = 1'h0;
    #10000;

    vif.RESETN         = 1'h1;
    #1000;
    wait(top_hdl.u_dut.sdr_init_done == 1);
    #1000;
    `uvm_info("DRV", "RESET applied", UVM_LOW)
  endtask

  // Task for the burst write operation.
  virtual task burst_write(sdram_item f_item);
    int i;
    $display("Start of burst_write task");
    @ (negedge vif.sys_clk);
    for (i = 0; i < f_item.bl; i++) begin
      vif.wb_stb_i = 1;
      vif.wb_cyc_i = 1;
      vif.wb_we_i = 1;
      vif.wb_sel_i = 4'b1111;
      vif.wb_addr_i = {f_item.Address[31:2] + i, 2'b00};
      $display("Bus signals activated.");

      vif.wb_dat_i = f_item.writte;
      f_item.writte += 100; 
      do begin
        @(posedge vif.sys_clk);
      end while (vif.wb_ack_o == 1'b0);
      @(negedge vif.sys_clk);
      $display("Burst number: %d, Write address: %h, Data written: %h", i, vif.wb_addr_i, vif.wb_dat_i);
    end
    vif.wb_stb_i = 0;
    vif.wb_cyc_i = 0;
    vif.wb_we_i = 'hx;
    vif.wb_sel_i = 'hx;
    vif.wb_addr_i = 'hx;
    vif.wb_dat_i = 'hx;
    $display("End of burst write process.");
  endtask

  // Task for the burst read operation.
  virtual task burst_read(bit[31:0] address);
    int j;
    $display("Start of burst_read task.");

    for (j = 0; j < 16; j++) begin
      vif.wb_stb_i = 1;
      vif.wb_cyc_i = 1;
      vif.wb_we_i = 0;
      vif.wb_addr_i = address + (j * 4);
      $display("Bus signals activated.");

      do begin
        @ (posedge vif.sys_clk);
      end while (vif.wb_ack_o == 1'b0);
      $display("Burst number: %d, ACK received for address %h, Data received: %h", j, vif.wb_addr_i, vif.wb_dat_o);
      @(negedge vif.sdram_clk);
    end
    vif.wb_stb_i = 0;
    vif.wb_cyc_i = 0;
    vif.wb_we_i = 'hx;
    vif.wb_addr_i = 'hx;
    $display("End of burst read process.");
  endtask
  
  // Task to print the contents of the memory.
  virtual task print_memory_contents();
    int address;
    int num_addresses = 1024;
    $display("Start of print_memory_contents task.");

    for (address = 0; address < num_addresses * 4; address += 4) begin
      vif.wb_stb_i = 1;
      vif.wb_cyc_i = 1;
      vif.wb_we_i = 0;
      vif.wb_addr_i = address;

      do begin
        @ (posedge vif.sys_clk);
      end while (vif.wb_ack_o == 1'b0);

      $display("Address: %h, Data read: %h", address, vif.wb_dat_o);
      @(negedge vif.sdram_clk);
    end

    vif.wb_stb_i = 0;
    vif.wb_cyc_i = 0;
    vif.wb_we_i = 'hx;
    vif.wb_addr_i = 'hx;

    $display("End of memory content read process.");
  endtask
endclass
